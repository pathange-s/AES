`timescale 1ns / 1ps

module sbox(inputByte, substitutedByte);
    
	input  [7:0] inputByte;
	output [7:0] substitutedByte;
    
	reg [7:0] substitutedByte;
    
    
    always @(inputByte)
    case (inputByte)
      8'h00: substitutedByte =8'h63;
	   8'h01: substitutedByte=8'h7c;
	   8'h02: substitutedByte=8'h77;
	   8'h03: substitutedByte=8'h7b;
	   8'h04: substitutedByte=8'hf2;
	   8'h05: substitutedByte=8'h6b;
	   8'h06: substitutedByte=8'h6f;
	   8'h07: substitutedByte=8'hc5;
	   8'h08: substitutedByte=8'h30;
	   8'h09: substitutedByte=8'h01;
	   8'h0a: substitutedByte=8'h67;
	   8'h0b: substitutedByte=8'h2b;
	   8'h0c: substitutedByte=8'hfe;
	   8'h0d: substitutedByte=8'hd7;
	   8'h0e: substitutedByte=8'hab;
	   8'h0f: substitutedByte=8'h76;
	   8'h10: substitutedByte=8'hca;
	   8'h11: substitutedByte=8'h82;
	   8'h12: substitutedByte=8'hc9;
	   8'h13: substitutedByte=8'h7d;
	   8'h14: substitutedByte=8'hfa;
	   8'h15: substitutedByte=8'h59;
	   8'h16: substitutedByte=8'h47;
	   8'h17: substitutedByte=8'hf0;
	   8'h18: substitutedByte=8'had;
	   8'h19: substitutedByte=8'hd4;
	   8'h1a: substitutedByte=8'ha2;
	   8'h1b: substitutedByte=8'haf;
	   8'h1c: substitutedByte=8'h9c;
	   8'h1d: substitutedByte=8'ha4;
	   8'h1e: substitutedByte=8'h72;
	   8'h1f: substitutedByte=8'hc0;
	   8'h20: substitutedByte=8'hb7;
	   8'h21: substitutedByte=8'hfd;
	   8'h22: substitutedByte=8'h93;
	   8'h23: substitutedByte=8'h26;
	   8'h24: substitutedByte=8'h36;
	   8'h25: substitutedByte=8'h3f;
	   8'h26: substitutedByte=8'hf7;
	   8'h27: substitutedByte=8'hcc;
	   8'h28: substitutedByte=8'h34;
	   8'h29: substitutedByte=8'ha5;
	   8'h2a: substitutedByte=8'he5;
	   8'h2b: substitutedByte=8'hf1;
	   8'h2c: substitutedByte=8'h71;
	   8'h2d: substitutedByte=8'hd8;
	   8'h2e: substitutedByte=8'h31;
	   8'h2f: substitutedByte=8'h15;
	   8'h30: substitutedByte=8'h04;
	   8'h31: substitutedByte=8'hc7;
	   8'h32: substitutedByte=8'h23;
	   8'h33: substitutedByte=8'hc3;
	   8'h34: substitutedByte=8'h18;
	   8'h35: substitutedByte=8'h96;
	   8'h36: substitutedByte=8'h05;
	   8'h37: substitutedByte=8'h9a;
	   8'h38: substitutedByte=8'h07;
	   8'h39: substitutedByte=8'h12;
	   8'h3a: substitutedByte=8'h80;
	   8'h3b: substitutedByte=8'he2;
	   8'h3c: substitutedByte=8'heb;
	   8'h3d: substitutedByte=8'h27;
	   8'h3e: substitutedByte=8'hb2;
	   8'h3f: substitutedByte=8'h75;
	   8'h40: substitutedByte=8'h09;
	   8'h41: substitutedByte=8'h83;
	   8'h42: substitutedByte=8'h2c;
	   8'h43: substitutedByte=8'h1a;
	   8'h44: substitutedByte=8'h1b;
	   8'h45: substitutedByte=8'h6e;
	   8'h46: substitutedByte=8'h5a;
	   8'h47: substitutedByte=8'ha0;
	   8'h48: substitutedByte=8'h52;
	   8'h49: substitutedByte=8'h3b;
	   8'h4a: substitutedByte=8'hd6;
	   8'h4b: substitutedByte=8'hb3;
	   8'h4c: substitutedByte=8'h29;
	   8'h4d: substitutedByte=8'he3;
	   8'h4e: substitutedByte=8'h2f;
	   8'h4f: substitutedByte=8'h84;
	   8'h50: substitutedByte=8'h53;
	   8'h51: substitutedByte=8'hd1;
	   8'h52: substitutedByte=8'h00;
	   8'h53: substitutedByte=8'hed;
	   8'h54: substitutedByte=8'h20;
	   8'h55: substitutedByte=8'hfc;
	   8'h56: substitutedByte=8'hb1;
	   8'h57: substitutedByte=8'h5b;
	   8'h58: substitutedByte=8'h6a;
	   8'h59: substitutedByte=8'hcb;
	   8'h5a: substitutedByte=8'hbe;
	   8'h5b: substitutedByte=8'h39;
	   8'h5c: substitutedByte=8'h4a;
	   8'h5d: substitutedByte=8'h4c;
	   8'h5e: substitutedByte=8'h58;
	   8'h5f: substitutedByte=8'hcf;
	   8'h60: substitutedByte=8'hd0;
	   8'h61: substitutedByte=8'hef;
	   8'h62: substitutedByte=8'haa;
	   8'h63: substitutedByte=8'hfb;
	   8'h64: substitutedByte=8'h43;
	   8'h65: substitutedByte=8'h4d;
	   8'h66: substitutedByte=8'h33;
	   8'h67: substitutedByte=8'h85;
	   8'h68: substitutedByte=8'h45;
	   8'h69: substitutedByte=8'hf9;
	   8'h6a: substitutedByte=8'h02;
	   8'h6b: substitutedByte=8'h7f;
	   8'h6c: substitutedByte=8'h50;
	   8'h6d: substitutedByte=8'h3c;
	   8'h6e: substitutedByte=8'h9f;
	   8'h6f: substitutedByte=8'ha8;
	   8'h70: substitutedByte=8'h51;
	   8'h71: substitutedByte=8'ha3;
	   8'h72: substitutedByte=8'h40;
	   8'h73: substitutedByte=8'h8f;
	   8'h74: substitutedByte=8'h92;
	   8'h75: substitutedByte=8'h9d;
	   8'h76: substitutedByte=8'h38;
	   8'h77: substitutedByte=8'hf5;
	   8'h78: substitutedByte=8'hbc;
	   8'h79: substitutedByte=8'hb6;
	   8'h7a: substitutedByte=8'hda;
	   8'h7b: substitutedByte=8'h21;
	   8'h7c: substitutedByte=8'h10;
	   8'h7d: substitutedByte=8'hff;
	   8'h7e: substitutedByte=8'hf3;
	   8'h7f: substitutedByte=8'hd2;
	   8'h80: substitutedByte=8'hcd;
	   8'h81: substitutedByte=8'h0c;
	   8'h82: substitutedByte=8'h13;
	   8'h83: substitutedByte=8'hec;
	   8'h84: substitutedByte=8'h5f;
	   8'h85: substitutedByte=8'h97;
	   8'h86: substitutedByte=8'h44;
	   8'h87: substitutedByte=8'h17;
	   8'h88: substitutedByte=8'hc4;
	   8'h89: substitutedByte=8'ha7;
	   8'h8a: substitutedByte=8'h7e;
	   8'h8b: substitutedByte=8'h3d;
	   8'h8c: substitutedByte=8'h64;
	   8'h8d: substitutedByte=8'h5d;
	   8'h8e: substitutedByte=8'h19;
	   8'h8f: substitutedByte=8'h73;
	   8'h90: substitutedByte=8'h60;
	   8'h91: substitutedByte=8'h81;
	   8'h92: substitutedByte=8'h4f;
	   8'h93: substitutedByte=8'hdc;
	   8'h94: substitutedByte=8'h22;
	   8'h95: substitutedByte=8'h2a;
	   8'h96: substitutedByte=8'h90;
	   8'h97: substitutedByte=8'h88;
	   8'h98: substitutedByte=8'h46;
	   8'h99: substitutedByte=8'hee;
	   8'h9a: substitutedByte=8'hb8;
	   8'h9b: substitutedByte=8'h14;
	   8'h9c: substitutedByte=8'hde;
	   8'h9d: substitutedByte=8'h5e;
	   8'h9e: substitutedByte=8'h0b;
	   8'h9f: substitutedByte=8'hdb;
	   8'ha0: substitutedByte=8'he0;
	   8'ha1: substitutedByte=8'h32;
	   8'ha2: substitutedByte=8'h3a;
	   8'ha3: substitutedByte=8'h0a;
	   8'ha4: substitutedByte=8'h49;
	   8'ha5: substitutedByte=8'h06;
	   8'ha6: substitutedByte=8'h24;
	   8'ha7: substitutedByte=8'h5c;
	   8'ha8: substitutedByte=8'hc2;
	   8'ha9: substitutedByte=8'hd3;
	   8'haa: substitutedByte=8'hac;
	   8'hab: substitutedByte=8'h62;
	   8'hac: substitutedByte=8'h91;
	   8'had: substitutedByte=8'h95;
	   8'hae: substitutedByte=8'he4;
	   8'haf: substitutedByte=8'h79;
	   8'hb0: substitutedByte=8'he7;
	   8'hb1: substitutedByte=8'hc8;
	   8'hb2: substitutedByte=8'h37;
	   8'hb3: substitutedByte=8'h6d;
	   8'hb4: substitutedByte=8'h8d;
	   8'hb5: substitutedByte=8'hd5;
	   8'hb6: substitutedByte=8'h4e;
	   8'hb7: substitutedByte=8'ha9;
	   8'hb8: substitutedByte=8'h6c;
	   8'hb9: substitutedByte=8'h56;
	   8'hba: substitutedByte=8'hf4;
	   8'hbb: substitutedByte=8'hea;
	   8'hbc: substitutedByte=8'h65;
	   8'hbd: substitutedByte=8'h7a;
	   8'hbe: substitutedByte=8'hae;
	   8'hbf: substitutedByte=8'h08;
	   8'hc0: substitutedByte=8'hba;
	   8'hc1: substitutedByte=8'h78;
	   8'hc2: substitutedByte=8'h25;
	   8'hc3: substitutedByte=8'h2e;
	   8'hc4: substitutedByte=8'h1c;
	   8'hc5: substitutedByte=8'ha6;
	   8'hc6: substitutedByte=8'hb4;
	   8'hc7: substitutedByte=8'hc6;
	   8'hc8: substitutedByte=8'he8;
	   8'hc9: substitutedByte=8'hdd;
	   8'hca: substitutedByte=8'h74;
	   8'hcb: substitutedByte=8'h1f;
	   8'hcc: substitutedByte=8'h4b;
	   8'hcd: substitutedByte=8'hbd;
	   8'hce: substitutedByte=8'h8b;
	   8'hcf: substitutedByte=8'h8a;
	   8'hd0: substitutedByte=8'h70;
	   8'hd1: substitutedByte=8'h3e;
	   8'hd2: substitutedByte=8'hb5;
	   8'hd3: substitutedByte=8'h66;
	   8'hd4: substitutedByte=8'h48;
	   8'hd5: substitutedByte=8'h03;
	   8'hd6: substitutedByte=8'hf6;
	   8'hd7: substitutedByte=8'h0e;
	   8'hd8: substitutedByte=8'h61;
	   8'hd9: substitutedByte=8'h35;
	   8'hda: substitutedByte=8'h57;
	   8'hdb: substitutedByte=8'hb9;
	   8'hdc: substitutedByte=8'h86;
	   8'hdd: substitutedByte=8'hc1;
	   8'hde: substitutedByte=8'h1d;
	   8'hdf: substitutedByte=8'h9e;
	   8'he0: substitutedByte=8'he1;
	   8'he1: substitutedByte=8'hf8;
	   8'he2: substitutedByte=8'h98;
	   8'he3: substitutedByte=8'h11;
	   8'he4: substitutedByte=8'h69;
	   8'he5: substitutedByte=8'hd9;
	   8'he6: substitutedByte=8'h8e;
	   8'he7: substitutedByte=8'h94;
	   8'he8: substitutedByte=8'h9b;
	   8'he9: substitutedByte=8'h1e;
	   8'hea: substitutedByte=8'h87;
	   8'heb: substitutedByte=8'he9;
	   8'hec: substitutedByte=8'hce;
	   8'hed: substitutedByte=8'h55;
	   8'hee: substitutedByte=8'h28;
	   8'hef: substitutedByte=8'hdf;
	   8'hf0: substitutedByte=8'h8c;
	   8'hf1: substitutedByte=8'ha1;
	   8'hf2: substitutedByte=8'h89;
	   8'hf3: substitutedByte=8'h0d;
	   8'hf4: substitutedByte=8'hbf;
	   8'hf5: substitutedByte=8'he6;
	   8'hf6: substitutedByte=8'h42;
	   8'hf7: substitutedByte=8'h68;
	   8'hf8: substitutedByte=8'h41;
	   8'hf9: substitutedByte=8'h99;
	   8'hfa: substitutedByte=8'h2d;
	   8'hfb: substitutedByte=8'h0f;
	   8'hfc: substitutedByte=8'hb0;
	   8'hfd: substitutedByte=8'h54;
	   8'hfe: substitutedByte=8'hbb;
	   8'hff: substitutedByte=8'h16;
	endcase
endmodule